module baugh_multi(a,b,p);   
